module my_dmux4way(b, c, d, e, a, sel[1:0]);
   input a;
   input [1:0] sel;

   output      b;
   output      c;
   output      d;
   output      e;

   // implementation

endmodule
