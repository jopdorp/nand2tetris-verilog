module my_dmux(a, b, i, s);
   input i, s;
   output a, b;

   // implementation

endmodule
