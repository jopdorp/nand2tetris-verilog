`ifndef half_adder
  `include "half_adder.sv"
`endif
`define full_adder 1

module full_adder(
    input  a,
    input  b,
    input  c,
    output carry,
    output sum
);

    // Put your code here

endmodule
