module or(c, a, b);
   input a, b;
   output c;

   // implementation

endmodule
