module not_n2t(output out, input in);
    nand gate1(out, in, in);
endmodule
