module dmux_8_way(
    input  in,
    input[2:0] sel,
    output[7:0] out
);

    // implementation

endmodule
