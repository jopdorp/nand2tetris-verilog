module my_and16(c[15:0], b[15:0], a[15:0]);
   input [15:0] a;
   input [15:0] b;
   output [15:0] c;
   
   // implementation

endmodule
