module my_not(b, a);
   input a;
   output b;

   // implementation
   
endmodule
