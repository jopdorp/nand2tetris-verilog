module test_alu();
   reg zx, zy, nx, ny, f, no;
   reg [15:0] x;
   reg [15:0] y;
   reg [15:0] exp_out;

   wire [15:0] out;
   
   alu u1(out, x, y, zx, zy, nx, ny, f, no);
   
   initial
     begin
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 1;
	nx = 0;
	zy = 1;
	ny = 0;
	f = 1;
	no = 0;
	exp_out = 16'b0000000000000000;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 1;
	nx = 1;
	zy = 1;
	ny = 1;
	f = 1;
	no = 1;
	exp_out = 16'b0000000000000001;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 1;
	nx = 1;
	zy = 1;
	ny = 0;
	f = 1;
	no = 0;
	exp_out = 16'b1111111111111111;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 0;
	nx = 0;
	zy = 1;
	ny = 1;
	f = 0;
	no = 0;
	exp_out = 16'b0000000000000000;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 1;
	nx = 1;
	zy = 0;
	ny = 0;
	f = 0;
	no = 0;
	exp_out = 16'b1111111111111111;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 0;
	nx = 0;
	zy = 1;
	ny = 1;
	f = 0;
	no = 1;
	exp_out = 16'b1111111111111111;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 1;
	nx = 1;
	zy = 0;
	ny = 0;
	f = 0;
	no = 1;
	exp_out = 16'b0000000000000000;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 0;
	nx = 0;
	zy = 1;
	ny = 1;
	f = 1;
	no = 1;
	exp_out = 16'b0000000000000000;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 1;
	nx = 1;
	zy = 0;
	ny = 0;
	f = 1;
	no = 1;
	exp_out = 16'b0000000000000001;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 0;
	nx = 1;
	zy = 1;
	ny = 1;
	f = 1;
	no = 1;
	exp_out = 16'b0000000000000001;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 1;
	nx = 1;
	zy = 0;
	ny = 1;
	f = 1;
	no = 1;
	exp_out = 16'b0000000000000000;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 0;
	nx = 0;
	zy = 1;
	ny = 1;
	f = 1;
	no = 0;
	exp_out = 16'b1111111111111111;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 1;
	nx = 1;
	zy = 0;
	ny = 0;
	f = 1;
	no = 0;
	exp_out = 16'b1111111111111110;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 0;
	nx = 0;
	zy = 0;
	ny = 0;
	f = 1;
	no = 0;
	exp_out = 16'b1111111111111111;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 0;
	nx = 1;
	zy = 0;
	ny = 0;
	f = 1;
	no = 1;
	exp_out = 16'b0000000000000001;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 0;
	nx = 0;
	zy = 0;
	ny = 1;
	f = 1;
	no = 1;
	exp_out = 16'b1111111111111111;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 0;
	nx = 0;
	zy = 0;
	ny = 0;
	f = 0;
	no = 0;
	exp_out = 16'b0000000000000000;

	#10
	x = 16'b0000000000000000;
	y = 16'b1111111111111111;
	zx = 0;
	nx = 1;
	zy = 0;
	ny = 1;
	f = 0;
	no = 1;
	exp_out = 16'b1111111111111111;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 1;
	nx = 0;
	zy = 1;
	ny = 0;
	f = 1;
	no = 0;
	exp_out = 16'b0000000000000000;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 1;
	nx = 1;
	zy = 1;
	ny = 1;
	f = 1;
	no = 1;
	exp_out = 16'b0000000000000001;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 1;
	nx = 1;
	zy = 1;
	ny = 0;
	f = 1;
	no = 0;
	exp_out = 16'b1111111111111111;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 0;
	nx = 0;
	zy = 1;
	ny = 1;
	f = 0;
	no = 0;
	exp_out = 16'b0101101110100000;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 1;
	nx = 1;
	zy = 0;
	ny = 0;
	f = 0;
	no = 0;
	exp_out = 16'b0001111011010010;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 0;
	nx = 0;
	zy = 1;
	ny = 1;
	f = 0;
	no = 1;
	exp_out = 16'b1010010001011111;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 1;
	nx = 1;
	zy = 0;
	ny = 0;
	f = 0;
	no = 1;
	exp_out = 16'b1110000100101101;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 0;
	nx = 0;
	zy = 1;
	ny = 1;
	f = 1;
	no = 1;
	exp_out = 16'b1010010001100000;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 1;
	nx = 1;
	zy = 0;
	ny = 0;
	f = 1;
	no = 1;
	exp_out = 16'b1110000100101110;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 0;
	nx = 1;
	zy = 1;
	ny = 1;
	f = 1;
	no = 1;
	exp_out = 16'b0101101110100001;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 1;
	nx = 1;
	zy = 0;
	ny = 1;
	f = 1;
	no = 1;
	exp_out = 16'b0001111011010011;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 0;
	nx = 0;
	zy = 1;
	ny = 1;
	f = 1;
	no = 0;
	exp_out = 16'b0101101110011111;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 1;
	nx = 1;
	zy = 0;
	ny = 0;
	f = 1;
	no = 0;
	exp_out = 16'b0001111011010001;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 0;
	nx = 0;
	zy = 0;
	ny = 0;
	f = 1;
	no = 0;
	exp_out = 16'b0111101001110010;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 0;
	nx = 1;
	zy = 0;
	ny = 0;
	f = 1;
	no = 1;
	exp_out = 16'b0011110011001110;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 0;
	nx = 0;
	zy = 0;
	ny = 1;
	f = 1;
	no = 1;
	exp_out = 16'b1100001100110010;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 0;
	nx = 0;
	zy = 0;
	ny = 0;
	f = 0;
	no = 0;
	exp_out = 16'b0001101010000000;

	#10
	x = 16'b0101101110100000;
	y = 16'b0001111011010010;
	zx = 0;
	nx = 1;
	zy = 0;
	ny = 1;
	f = 0;
	no = 1;
	exp_out = 16'b0101111111110010;
     end

   initial
     $monitor("alu %d %b %b %b %b %b %b %b %b (%b %b)", $time, zx, zy, nx, ny, f, no, x, y, out, exp_out);
   
endmodule
