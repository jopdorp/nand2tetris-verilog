module not_n2t(input in, output out);
    nand not_n2t(out, in, in);
endmodule
