module my_and(c, a, b);
   input a, b;
   output c;

   // implementation

endmodule 
