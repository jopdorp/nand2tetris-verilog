module or_8_way(b, a[7:0]);
   input [7:0] a;
   output b;

   // implementation

endmodule
