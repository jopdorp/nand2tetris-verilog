module main;
   initial
     begin
	$display("whats up world");
	$finish ;
     end
endmodule
