module my_mux16(c[15:0], a[15:0], b[15:0], s);
   input [15:0] a;
   input [15:0] b;
   input 	s;
   output [15:0] c;

   // implementation

endmodule
