module add16(c, a, b);
   input [15:0] a;
   input [15:0] b;
   output [15:0] c;

   // Put your code here:

endmodule
