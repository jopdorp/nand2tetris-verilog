module not_16(b[15:0], out[15:0]);
   input [15:0] a;
   output [15:0] b;

endmodule
