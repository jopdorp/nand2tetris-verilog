module dmux_4_way(input in, input[1:0] sel, output[7:0] out);

   // implementation

endmodule
