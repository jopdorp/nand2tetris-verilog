module my_or(c, a, b);
   input a, b;
   output c;

   // implementation

endmodule
