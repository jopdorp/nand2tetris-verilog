module bit_n2t(in, load, reset, clk, out, );
   input in, load, clk, reset;
   output out;

endmodule
