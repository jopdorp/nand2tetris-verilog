module bit(out, in, load, reset, clk);
   input in, load, clk, reset;
   output out;

   // implementation

endmodule
