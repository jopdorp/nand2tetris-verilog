module my_or8way(b, a[7:0]);
   input [7:0] a;
   output b;

   // implementation

endmodule
