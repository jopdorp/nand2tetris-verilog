module xor_n2t(output out, input a, input b);

   // implementation

endmodule
