module dmux_8_way(b, c, d, e, f, g, h, j, a, sel[2:0]);
   input a;
   input [2:0] sel;

   // implementation

endmodule
