module not_n2t(input in, output out);
    nand result(out, in, in);
endmodule
