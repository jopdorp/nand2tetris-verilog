module dff(out, data, clk);
   input data, clk;
   output out;
   reg 	  out;

   // Put your code here:

endmodule
