//This file is here to verify that you installed and configured you environment correctly.
module hello_verilog_tb;

   initial begin
      $display("Hello world!");
   end

endmodule
