module my_mux(c, a, b, s);
   input a, b, s;
   output c;

   // implementation

endmodule
