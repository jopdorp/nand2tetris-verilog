module alu(out, zr, ng, x, y, zx, zy, nx, ny, f, no);
   input [15:0] x;
   input [15:0] y;
   input zx, zy, nx, ny, f, no;

   output [15:0] out;
   output 	 zr, ng;

   // implementation

endmodule
