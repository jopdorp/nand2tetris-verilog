module not_n2t(in, out);
    input in;
    input out;

    nand gate1(out, in, in);

endmodule
