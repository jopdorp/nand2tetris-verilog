module my_mux4way16(e[15:0], a[15:0], b[15:0], c[15:0], d[15:0], sel[1:0]);
   input [15:0] a;
   input [15:0] b;
   input [15:0] c;
   input [15:0] d;
   input [1:0] sel;

   output [15:0] e;

   // implementation

endmodule
