module inc16(b, a);
   input [15:0] a;
   output [15:0] b;

   // Put your code here:

endmodule
