module register(out, in, load, reset, clk);
   input [15:0] in;
   input load, clk, reset;
   output [15:0] out;

   // implementation

endmodule
