module and(c, a, b);
   input a, b;
   output c;

   // implementation

endmodule 
