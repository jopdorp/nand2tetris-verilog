module bit_n2t(out, in, load, reset, clk);
   input in, load, clk, reset;
   output out;

   // Put your code here:

endmodule
