module ram8(out, in, addr, load, clk);
   input [15:0] in;
   input [2:0] 	addr;
   input 	load, clk;
   output [15:0] out;

   // Put your code here:

endmodule
