module my_xor(c, a, b);
   input a, b;
   output c;

   // implementation

endmodule
