module half_adder(a, b, ca, s);
   input a, b;
   output ca, s;

   // Put your code here:

endmodule
