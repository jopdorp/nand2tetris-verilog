module full_adder(ca, s, a, b, c);
   input a, b, c;
   output ca, s;

   // implementation

endmodule
