module my_not16(b[15:0], a[15:0]);
   input [15:0] a;
   output [15:0] b;

   // implementation

endmodule
