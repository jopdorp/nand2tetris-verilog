module full_adder(ca, s, a, b, c);
   input a, b, c;
   output ca, s;

   // Put your code here:

endmodule
