`ifndef xor_n2t
  `include "../01/xor_n2t.sv"
`endif
`define half_adder 1

module half_adder(
    input  a,
    input  b,
    output carry,
    output sum
);

    // Put your code here

endmodule