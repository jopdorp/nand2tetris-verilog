module half_adder(a, b, ca, s);
   input a, b;
   output ca, s;

   // implementation

endmodule
